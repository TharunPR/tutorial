module counter(a,b,count);

endmodule